`include "para_defines.v"

module ysyx_23060124_lsu(
  input                               i_clk   ,
  input                               i_rst_n , 
  input [`ysyx_23060124_ISA_WIDTH - 1:0] lsu_src2,
  input [`ysyx_23060124_ISA_WIDTH - 1:0] alu_res,
  input [`ysyx_23060124_OPT_WIDTH - 1:0] load_opt,
  input [`ysyx_23060124_OPT_WIDTH - 1:0] store_opt,
  output reg [`ysyx_23060124_ISA_WIDTH - 1:0] lsu_res
);
reg [`ysyx_23060124_ISA_WIDTH - 1:0] read_res, store_res;

//   wire ren = |load_opt;
//   wire [`ysyx_23060124_OPT_WIDTH-1:0] raddr = alu_res;
//   wire [32-1:0] rdata;
//   always @(*) begin
//     case (load_opt)
//       `ysyx_23060124_OPT_LSU_LB:  lsu_res = {{24{rdata[ 7]}}, rdata[ 7:0]};
//       `ysyx_23060124_OPT_LSU_LH:  lsu_res = {{16{rdata[15]}}, rdata[15:0]};
//       `ysyx_23060124_OPT_LSU_LW:  lsu_res = rdata;
//       `ysyx_23060124_OPT_LSU_LBU: lsu_res = {24'b0, rdata[ 7:0]};
//       `ysyx_23060124_OPT_LSU_LHU: lsu_res = {16'b0, rdata[15:0]};
//       default:  lsu_res = `ysyx_23060124_OPT_WIDTH'b0;
//     endcase
//   end

//   reg  [7:0] mask;
//   wire [7:0] wmask;
//   wire [32-1:0] waddr,wdata;
//   always @(*) begin
//     case (store_opt)
//       `ysyx_23060124_OPT_LSU_SB:  mask = 8'b0000_0001;
//       `ysyx_23060124_OPT_LSU_SH:  mask = 8'b0000_0011;
//       `ysyx_23060124_OPT_LSU_SW:  mask = 8'b0000_1111;
//       default:  mask = 8'b0;
//     endcase
//   end

import "DPI-C" function void npc_pmem_read (input int raddr, output int rdata, input bit ren, input int len);
import "DPI-C" function void npc_pmem_write (input int waddr, input int wdata, input bit wen, input int len);
//   always @(*) begin
//     npc_pmem_write(waddr, wdata, 1, wmask);
//     npc_pmem_read (raddr, rdata, ren, 4);
//   end
//store

// always @(alu_res) begin
//     case(store_opt)
//     `ysyx_23060124_OPT_LSU_SB: begin store_res={24'b0, lsu_src2[7:0]}; end
//     `ysyx_23060124_OPT_LSU_SH: begin store_res={16'b0, lsu_src2[15:0]}; end
//     `ysyx_23060124_OPT_LSU_SW: begin store_res=lsu_src2; end
//     endcase
// end
reg [`ysyx_23060124_ISA_WIDTH - 1 : 0] store_addr, store_src2;
reg [`ysyx_23060124_OPT_WIDTH - 1 : 0] store_opt_next;

//load
// always @(alu_res) begin
//     case(load_opt)
//     `ysyx_23060124_OPT_LSU_LB: begin  npc_pmem_read(alu_res, read_res, |load_opt, 1); end
//     `ysyx_23060124_OPT_LSU_LH: begin  npc_pmem_read(alu_res, read_res, |load_opt, 2); end
//     `ysyx_23060124_OPT_LSU_LW: begin  npc_pmem_read(alu_res, read_res, |load_opt, 4); end
//     `ysyx_23060124_OPT_LSU_LBU: begin  npc_pmem_read(alu_res, read_res, |load_opt, 1); end
//     `ysyx_23060124_OPT_LSU_LHU: begin  npc_pmem_read(alu_res, read_res, |load_opt, 2); end
//     default: begin read_res = `ysyx_23060124_ISA_WIDTH'b0; end
//     endcase
// end

always @(*) begin
    case(load_opt)
    `ysyx_23060124_OPT_LSU_LB: begin lsu_res = {{24{read_res[7]}}, read_res[7:0]}; end
    `ysyx_23060124_OPT_LSU_LH: begin lsu_res = {{16{read_res[15]}}, read_res[15:0]}; end
    `ysyx_23060124_OPT_LSU_LW: begin lsu_res =read_res; end
    `ysyx_23060124_OPT_LSU_LBU: begin lsu_res = {24'b0, read_res[7:0]}; end
    `ysyx_23060124_OPT_LSU_LHU: begin lsu_res = {{16'b0}, read_res[15:0]}; end
    default: begin lsu_res = `ysyx_23060124_ISA_WIDTH'b0; end
    endcase
end

ysyx_23060124_Reg #(`ysyx_23060124_ISA_WIDTH + `ysyx_23060124_ISA_WIDTH + `ysyx_23060124_OPT_WIDTH,  0) lsu_reg(
  .clk(i_clk),
  .rst(i_rst_n),
  .din({alu_res, store_opt, lsu_src2}),
  .dout({store_addr,store_opt_next, store_src2}),
  .wen(1)
);

always @(*) begin
    case(store_opt_next)
    `ysyx_23060124_OPT_LSU_SB: begin  npc_pmem_write(store_addr, store_src2, |store_opt_next, 1); end
    `ysyx_23060124_OPT_LSU_SH: begin  npc_pmem_write(store_addr, store_src2, |store_opt_next, 2); end
    `ysyx_23060124_OPT_LSU_SW: begin  npc_pmem_write(store_addr, store_src2, |store_opt_next, 4); end
    endcase
end

always @(*) begin
  npc_pmem_read(alu_res, read_res, |load_opt, 4);
end

endmodule
