module ysyx_23060124_AGU (
    input              [32-1:0]         src1                       ,
    input              [32-1:0]         src2                       ,
    output             [32-1:0]         res                         
);

assign res =  src1 + src2;

endmodule
